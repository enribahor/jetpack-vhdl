------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : barryair.ppm 
--- Filas    : 32 
--- Columnas : 16 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_barryair is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(9-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_barryair;


architecture BEHAVIORAL of ROM_RGB_9b_barryair is
  signal addr_int  : natural range 0 to 2**9-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "011010001",
       "110101010",
       "011010001",
       "111111111",
       "111111111",
       "011010001",
       "011010001",
       "001000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "011010001",
       "111111101",
       "110101010",
       "011010001",
       "111111111",
       "001000000",
       "011010001",
       "001000000",
       "011010001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "001000000",
       "110101010",
       "110101010",
       "110101010",
       "110101010",
       "011010001",
       "011010001",
       "011010001",
       "011010001",
       "001000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "011010001",
       "011010001",
       "110101010",
       "110101010",
       "001000000",
       "011010001",
       "001000000",
       "001000000",
       "001000000",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "011010001",
       "110101010",
       "110101010",
       "110101010",
       "001000000",
       "011010001",
       "001000000",
       "001000000",
       "011010001",
       "100100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "011010001",
       "011010001",
       "011010001",
       "011010001",
       "011010001",
       "001000000",
       "001000000",
       "001000000",
       "110101101",
       "111111101",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "001000000",
       "110101010",
       "011010001",
       "011010001",
       "011010001",
       "001000000",
       "001000000",
       "001000000",
       "110101101",
       "011010001",
       "011010001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "001000000",
       "110101010",
       "011010001",
       "011010001",
       "011010001",
       "001000000",
       "001000000",
       "001000000",
       "111111101",
       "001000000",
       "011010001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "001000000",
       "110101010",
       "100100011",
       "110101010",
       "100100011",
       "001000000",
       "001000000",
       "001000000",
       "111111101",
       "011010001",
       "001000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "001000000",
       "110101010",
       "100100011",
       "110101010",
       "010010010",
       "000000000",
       "110101101",
       "001000000",
       "111111101",
       "111111101",
       "001000000",
       "111111101",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "001000000",
       "110101010",
       "100100011",
       "110101010",
       "010010010",
       "001000000",
       "111111101",
       "011010001",
       "111111101",
       "111111101",
       "111111101",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "011010001",
       "011010001",
       "100100011",
       "010010010",
       "010010010",
       "001000000",
       "111111101",
       "111111101",
       "111111101",
       "111111101",
       "111111101",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "011010001",
       "011010001",
       "100100011",
       "100100011",
       "100100011",
       "001000000",
       "001000000",
       "111111101",
       "111111101",
       "111111101",
       "011010001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "001000000",
       "011010001",
       "100100011",
       "100100011",
       "100100011",
       "001000000",
       "001000000",
       "001000000",
       "100100011",
       "000000000",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "011010001",
       "100100011",
       "100100011",
       "100100011",
       "000000000",
       "110101101",
       "111111101",
       "001000000",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100011",
       "000000000",
       "100100011",
       "100100011",
       "000000000",
       "111111101",
       "111111101",
       "100100011",
       "100100011",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "000000000",
       "100100011",
       "100100011",
       "001000000",
       "111111101",
       "111111101",
       "111111101",
       "111111101",
       "111111101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "000000000",
       "011010001",
       "110101101",
       "000000000",
       "110101101",
       "110101101",
       "110101101",
       "110101101",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "000000000",
       "001000000",
       "001000000",
       "010010010",
       "000000000",
       "011010001",
       "100100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "001000000",
       "001000000",
       "000000000",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "001000000",
       "001000000",
       "000000000",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "000000000",
       "111111111",
       "000000000",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "001000000",
       "111111111",
       "000000000",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "010010010",
       "000000000",
       "111111111",
       "000000000",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010010010",
       "000000000",
       "111111111",
       "111111111",
       "000000000",
       "100100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100011",
       "010010010",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

