------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : nivelfuegoBW.ppm 
--- Filas    : 256 
--- Columnas : 1024 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_nivelfuegoBW is
  port (
    clk  				: in  std_logic;   -- reloj
	 bloquea				  : in std_logic; 	--se�al que indica si se bloquean las primeras 256 posiciones
    addr, addr_munyeco  : in  std_logic_vector(18-1 downto 0);
    dout, dout_munyeco  : out std_logic 
  );
end ROM_RGB_9b_nivelfuegoBW;


architecture BEHAVIORAL of ROM_RGB_9b_nivelfuegoBW is
  signal addr_int, addr_munyeco_int  : natural range 0 to 2**18-1;
	signal rango : std_logic_vector(9 downto 0);
	signal rango_munyeco : std_logic_vector(9 downto 0);
	signal rango_int : natural range 0 to 2**12-1;
	signal rango_int_munyeco : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic;
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '1',
       '1',
       '1',
       '1',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0',
       '0'
        );

begin



  addr_int <= TO_INTEGER(unsigned(addr));
  addr_munyeco_int <= TO_INTEGER(unsigned(addr_munyeco));
 -- bloquea_avanza <= addr - "00000000"&avanza_obstaculo;
	--bloquea_int <= TO_INTEGER(unsigned(bloquea_avanza));
	rango <= addr(9 downto 0);
	rango_int <= TO_INTEGER(unsigned(rango));
	rango_munyeco <= addr_munyeco(9 downto 0);
	rango_int_munyeco <= TO_INTEGER(unsigned(rango_munyeco));
  P_ROM: process (clk)
  begin
	 if clk'event and clk='1' then
		if bloquea = '1' then
			--if addr(9 downto 8) = "00" then
			if rango_int < 512 then
				dout <= '0';
			else 
				dout <= filaimg(addr_int);
			end if;
			if rango_int_munyeco < 512 then
				dout_munyeco <= '0';
			else dout_munyeco <= filaimg(addr_munyeco_int);
			end if;
			--if addr_munyeco(9 downto 8) = "00" then
			--if addr_munyeco(9 downto 0) < "0100000000" then
			--	dout_munyeco <= '0';
			--else dout_munyeco <= filaimg(addr_munyeco_int);
			--end if;
		else
			dout <= filaimg(addr_int);
			dout_munyeco <= filaimg(addr_munyeco_int);
		end if;
		--dout <= '0';
		--dout_munyeco <= '0';
	 end if;
  end process;
end BEHAVIORAL;



--
--  addr_int <= TO_INTEGER(unsigned(addr));
--  addr_munyeco_int <= TO_INTEGER(unsigned(addr_munyeco));
--
--  P_ROM: process (clk)
--  begin
--	 if clk'event and clk='1' then
--		if bloquea = '1' then
--			if addr(9 downto 8) = "00" then
--				dout <= '0';
--			else dout <= filaimg(addr_int);
--			end if;
--			--if addr_munyeco(9 downto 8) = "00" then
--			if addr_munyeco(9 downto 0) < "0100000000" then
--				dout_munyeco <= '0';
--			else dout_munyeco <= filaimg(addr_munyeco_int);
--			end if;
--		else
--			dout <= filaimg(addr_int);
--			dout_munyeco <= filaimg(addr_munyeco_int);
--		end if;
--		--dout <= '0';
--		--dout_munyeco <= '0';
--	 end if;
--  end process;


